module AGU (
    input [15:0] H0, // Horizontal offset
    input [15:0] V0, // Vertical offset
    input [15:0] SW, // Source Width
    input [15:0] SH, // Source Height
    input [15:0] TW, // Target Width
    input [15:0] TH, // Target Height
    output [13:0] SRAM_addr, // Address to SRAM
);





endmodule